`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Boston University
// Engineer: Jackson Clary
// 
// Create Date: 10/01/2024 02:20:25 PM
// Design Name: Carry-Select-Adder
// Module Name: CSA_64bit_tb_0
// Project Name: EC413 Lab 3
//////////////////////////////////////////////////////////////////////////////////


module CSA_64bit_tb_0;

    reg [63:0] a, b;
    reg c_in;
    
    wire [63:0] sum;
    wire c_out;
    
    CSA2_64bit_0 uut (
        .a(a),
        .b(b),
        .c_in(c_in),
        .sum(sum),
        .c_out(c_out)
    );
    
    integer i;
    initial begin
        
        a = 64'h0000000000000003;
        b = 64'h0000000000000005;
        c_in = 0;
        #10;
        
        a = 64'h0000000000000003;
        b = 64'h0000000000000005;
        c_in = 1;
        #10;
        
        a = 64'hFFFFFFFFFFFFFFFF;
        b = 64'h0000000000000001;
        c_in = 1;
        #10;
        
        a = 64'h000000000000000A;
        b = 64'hFFFFFFFFFFFFFFF6;
        c_in = 0;
        #10;
        
        a = 64'hFFFFFFFFFFFFFFFF;
        b = 64'hFFFFFFFFFFFFFFFF;
        c_in = 1;
        #10;
        
        a = 64'b0;
        b = 64'b0;
        c_in = 1'b0;
        

        for (i = 0; i < 12; i = i +1) begin
            a = $random;
            b = $random;
            c_in = $random % 2;
            #10;
        end
        $finish;
    end
endmodule
